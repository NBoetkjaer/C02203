-- -----------------------------------------------------------------------------
--
--  Title      : Finite state machine and datapath of the GCD
--             :
--  Developers : Anders Greve(s073188) and Nicolas B�tkj�r (s918819) 
-- 		      :
--  Purpose    : This design is the FSM and Datapath of the Greatest Common Divisor
--             :
--  Notes      : Implementation of Euclids GCD algorithm with repeated subtration.
--             : The implementation is speed optimized, by using a Mealy state (CmpAB)
--             : and thereby removing states in inner 'loop' of the algorithm.
--             :
--  Revision   :  02203 fall 2014 v.1
--              
-- -----------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY gcd IS            
    PORT (clk:      IN std_logic;				-- The clock signal.
          reset:    IN std_logic;				-- Reset the module.
          req:      IN std_logic;				-- Start computation.
          AB:       IN unsigned(7 downto 0);	-- The two operands.
          ack:      OUT std_logic;				-- Computation is complete.
          C:        OUT unsigned(7 downto 0));	-- The result.  
END gcd;

architecture FSMD_optim of gcd is
-- FSMD States 
type state_type is ( InputA, LoadA, RegAdone, InputB, LoadB, CmpAB, DoneC );
-- Declare signals
signal reg_a,next_reg_a,next_reg_b,reg_b : unsigned(7 downto 0);
signal state, next_state : state_type; 
signal diff_ab, diff_ba : signed(8 downto 0); -- One extra bit to hold the sign-bit.

begin
	diff_ab <= signed(('0' & reg_a)) - signed(('0' & reg_b));
	diff_ba <= signed(('0' & reg_b)) - signed(('0' & reg_a));
	
	-- Combinatoriel logic
	CL: process (req, AB, state, reg_a, reg_b, diff_ab, diff_ba, reset)
	begin
		next_reg_a <= reg_a;
		next_reg_b <= reg_b;
		ack <= '0';	
		C <= (others =>'Z');		
		case (state) is
		
		When InputA =>
			if req = '1' then
				next_state <= LoadA;
			else
				next_state <= InputA;
			end if;
		  
		When LoadA =>  
			next_state <= RegAdone;
			next_reg_a <= AB;
			
		When RegAdone =>
			ack <= '1';
			if req = '0' then
				next_state <= InputB;
			else
				next_state <= RegAdone;
			end if;      
		
		When InputB =>
			if req = '1' then
				next_state <= LoadB;
			else
				next_state <= InputB;
			end if;     
		  
		When LoadB=>
			next_reg_b <= AB;
			next_state <= CmpAB;
		  
		When CmpAB =>
			if diff_ab(8) = '1' then -- If sign bit is set b > a
				next_reg_b <= unsigned(diff_ba(7 downto 0));
				next_state <= CmpAB;		
			elsif diff_ab(7 downto 0) = 0 then			
				next_state <= DoneC;
			else 
				next_reg_a <= unsigned(diff_ab(7 downto 0));
				next_state <= CmpAB;
			end if;
				
		When DoneC =>
			ack <= '1';
			C <= reg_a;
			if req = '0' then
				next_state <= InputA;
			else
				next_state <= DoneC;
			end if;  
			
	   end case;      
	end process CL; 

	-- Registers
	seq: process (clk, reset)
	begin
		if reset = '1' then
			state <= InputA;         -- Reset to initial state 
		elsif rising_edge(clk) then
			state <= next_state;
			reg_a <= next_reg_a;
			reg_b <= next_reg_b;
		end if;
	end process seq;
	
end FSMD_optim;

